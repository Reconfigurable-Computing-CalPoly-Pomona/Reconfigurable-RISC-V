`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/17/2019 04:19:47 PM
// Design Name: 
// Module Name: axi_pkg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// Contains the interface and types defined for the AXI 4 Protocol
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// TODO
module axi_pkg(

    );
endmodule
