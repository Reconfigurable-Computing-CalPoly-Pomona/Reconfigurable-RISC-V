//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Ben Kueffler
// 
// Create Date: 04/21/2019 11:37:42 AM
// Design Name: multicore
// Module Name: hazard_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description:
// Handles data, control, and structural hazards that occur as a part of the pipelining
// nature of the processor
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module hazard_unit(
  // System clock
  logic i_aclk,

  // Asynchronous reset
  logic i_areset_n
);
endmodule
